module controller(output );

endmodule
